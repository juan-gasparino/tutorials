//Tutorial_1

module hello_world();

  initial begin
    $display("\n\t testing\n");
  end

endmodule